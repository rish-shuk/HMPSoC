    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984�N`    ���    �y�X�[#)$]p(.ozb�2`�,AY&,9�~kFu�"*u�j��2cf%(F�H�q��S����7?�>��Ѳ����?���S�=L�,�	��

Y����     
������