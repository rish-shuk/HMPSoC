    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;1342179840�N`    ��    ��R5�P%�U [׌�jR����B=���"�q=���p��փ�n�#��@�Sɖ;��r�d�kE���n}/H����a�l
c��E��,

Y����     
�5����