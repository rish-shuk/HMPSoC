    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984��N`    U� 7    ��W��y�&�t���g�u��
���mLW����B��{�bC���M5`����0�VK&]*@�����f�3o�4���K��

Y����     
�6��̾