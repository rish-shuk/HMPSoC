    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984ހN`    %5+    �zץ�ƽ�Ѯ�(��&B2U��a��ǣ,O
%��W,Q�W��q�CA�S��l�卵��M;�g���cf��*SW�iPEsn2b�%!�X�_

Y����     
�����(