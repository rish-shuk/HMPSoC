    Mac OS X            	   2  I     {                                      ATTR      {  X  #                 X   �  "com.apple.LaunchServices.OpenWith      �     com.apple.TextEncoding     �     com.apple.lastuseddate#PS         Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     a     com.dropbox.attrs    bplist00�WversionTpath_bundleidentifier _!/System/Applications/TextEdit.app_com.apple.TextEdit/1U                            jutf-8;134217984T�f    nƍ    ����"3���l�a���ݤ�ӈ�� Vv�'6��x�1�^g)6��j�*w��BE��I4�x��R��I��� ��J[n�ڔ�����

Y����     
����Ӑ