    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984U�f    ��-    �}�ɐ�iD��y�(�)�Q�P��ۉ�&�Wޙ+����aq����L$ |�����7����t�0��W���2�������I�GB\

Y����     
�7θІ