    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984�N`    �IC4    �B�u�Qt��d�h�rjnaT���S0��������d�<�()yC����oC������,�^Ł��3C��kV��5r��

Y����     
�4����