package macros is
    constant data_width : integer := 12;
    constant sampling_rate : integer := 16000;
    constant sampling_delay : integer := 6249;
end package macros;