    Mac OS X            	   2  I     {                                      ATTR      {  X  #                 X   �  "com.apple.LaunchServices.OpenWith      �     com.apple.TextEncoding     �     com.apple.lastuseddate#PS         Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     a     com.dropbox.attrs    bplist00�WversionTpath_bundleidentifier _!/System/Applications/TextEdit.app_com.apple.TextEdit/1U                            jutf-8;134217984�f    9:�8    �D�s�R��E������<o:!�Pr���i�����x5NN�ӏL?@�u|��f9mc�%��}K}	���ȭ8�PV�1%Ȝ�+w�JD

Y����     
�:����