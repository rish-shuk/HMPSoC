    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   Y  7com.apple.metadata:kMDLabel_c6abldq2zv5c2u5ebywntxmkue     �     com.dropbox.attrs    utf-8;134217984؇f    �8    򴜜�T�v��ໜ7I�1(q`�`Y��`�Mu�"��A*}i:Lo�v���6����A�K����6]⪥'�A��U2�֚}N�^��

Y����     
�<Ƌ��