    Mac OS X            	   2   �                                           ATTR         �   9                  �     com.apple.TextEncoding      �     com.apple.lastuseddate#PS           com.dropbox.attrs    utf-8;134217984��f    H/"    

Y����     
�9�ⰻ